library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MIPS is
    Port (
		
	 );
end MIPS;

architecture rtl of MIPS is
begin
    
end rtl;